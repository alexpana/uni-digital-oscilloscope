--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   08:28:10 06/07/2013
-- Design Name:   
-- Module Name:   E:/SEM2/SSC/project-repo/uni-digital-oscilloscope/testproj/ttr/osc/testRandgen.vhd
-- Project Name:  osc
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: randgen
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY testRandgen IS
END testRandgen;
 
ARCHITECTURE behavior OF testRandgen IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT randgen
    PORT(
         startBit : IN  std_logic;
         reqBit : IN  std_logic;
         rbit : OUT  std_logic;
         rbitValid : OUT  std_logic;
         clk : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal startBit : std_logic := '0';
   signal reqBit : std_logic := '0';
   signal clk : std_logic := '0';

 	--Outputs
   signal rbit : std_logic;
   signal rbitValid : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: randgen PORT MAP (
          startBit => startBit,
          reqBit => reqBit,
          rbit => rbit,
          rbitValid => rbitValid,
          clk => clk
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;
		
		reqBit <= '1';
		wait for clk_period * 300;		
		reqBit <= '0';
		wait for clk_period * 300;		
		reqBit <= '1';
		wait for clk_period * 300;

      -- insert stimulus here 

      wait;
   end process;

END;
