library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity color_select is
	port (
		x, y:			in std_logic_vector(10 downto 0);
		sel:			out std_logic
	);
end color_select;

architecture Behavioral of color_select is

begin

	

end Behavioral;

